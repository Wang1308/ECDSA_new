import elliptic_curve_structs::*;

module point_add (
	input 	logic 			clk, Reset,
	//input  	curve_point_t 	P, Q,
	input 	logic [255:0]  	P_x,
	input 	logic [255:0]  	P_y,
	input 	logic [255:0]  	Q_x,
	input 	logic [255:0]  	Q_y,
	input   curve_parameters_t params,
	output 	logic 			Done,
	//output 	curve_point_t 	R
	output 	logic [255:0]  	R_x,
	output 	logic [255:0]  	R_y
);

	logic mult0_done, inv_done, mult1_done, mult2_done;
	logic[255:0] sum0, sum1, sum2, sum3, sum4, sum5, sum6, sum7, sum8, s;
	logic[255:0] inv1;
	logic[255:0] prod1, prod2, prod3;
	logic reset0, reset1, reset2, inv_reset;

	logic[2:0] counter;

	//s = (Py + Qy) / (Px + Qx)
	//Rx = s*s + s + Px + Qx
	//Ry = s(Px + Rx) + Rx + Py

	// s = (Py - Qy) / (Px - Qx)
	// Rx = s*s - Px - Qx
	// Ry = s(Px - Rx) - Py

	/* code for testbench */
	always_ff @ (posedge clk)
	begin
		if(Reset) begin
			counter <= 0;
			reset2 <= 1'b0;
		end

		else
		begin
			if(mult1_done)
				counter <= counter + 1'b1;
			if(counter > 5)
				reset2 <= 1'b1;
		end
	end

	add add0(.a(P_y), .b(Q_y), .params(params), .op(1'b1), .sum(sum0));	// Py - Qy
	add add1(.a(P_x), .b(Q_x), .params(params), .op(1'b1), .sum(sum1));	// Px - Qx
	modular_inverse inv0(.clk(clk), .Reset(Reset), .in( sum1), .params(params), .out(inv1), .Done(inv_done)); //1/Px-Qx

	multiplier mult0(.clk, .Reset(~inv_done | Reset), .a(sum0), .b(inv1), .params(params), .Done(mult0_done), .product(s)); //slope

	multiplier mult1(.clk, .Reset(~mult0_done | Reset), .a(s), .b(s), .params(params), .Done(mult1_done), .product(prod2)); // s^2
	add add2(.a(P_x), .b(Q_x), .params(params), .op(1'b0), .sum(sum3));	// Px + Qx
	add add3(.a(prod2), .b(sum3), .params(params), .op(1'b1), .sum(sum4)); // s^2 - (Px + Qx)
	add add4(.a(P_x), .b(sum4), .params(params), .op(1'b1), .sum(sum5));	// Px - Rx
	add add5(.a(prod3), .b(P_y), .params(params), .op(1'b1), .sum(sum6)); // s(Px-Rx) - Py
	multiplier mult2(.clk, .Reset(~reset2 | Reset), .a(s), .b(sum5), .params(params), .Done(mult2_done), .product(prod3)); //s(Px - Rx)
	/* to use a nonzero a, uncomment below line and replace all "sum4" with "sum8" */
	//add #(17) 
	add add7(.a(sum4), .b(params.p), .params(params), .op(1'b0/*1'b0*/), .sum(sum8)); // Rx + a (for x^3 + 2x + 2, a is 2) //


	assign R_x = sum8;
	assign R_y = sum6;
	assign Done = mult0_done & inv_done & mult1_done & mult2_done;

endmodule

